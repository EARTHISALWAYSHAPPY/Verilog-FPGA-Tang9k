//File name : 
//Description : 
//Company :
//Project :
//-------------------     |     NEW
//Version :               |
//Date :                  |
//Author :                |
//Remark :                |   
//-------------------     |   
//Version :               |
//Date :                  |
//Author :                |
//Remark :                |     OLD
                          V
module moduleName (
   
);
//-------------------  
// Constant Declaration 
// for initial Const.
//-------------------

//-------------------  
// Signal Declaration 
// for initial reg,wire
//-------------------

//-------------------  
// Output 
// assignd wire <= reg
//-------------------

//-------------------  
// Process Declaration
// @always
//-------------------
endmodule